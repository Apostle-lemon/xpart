`timescale 1ns / 1ps

module vga_gen_grafic(
        input               clk,
        input               rst_n,

        input [7:0] char_1,
        input [7:0] char_2,
        input [7:0] char_3,
        input [7:0] char_4,
        input [7:0] char_5,
        input [7:0] char_6,
        input [7:0] char_7,
        input [7:0] char_8,
        input [7:0] char_9,
        input [7:0] char_10,
        input [7:0] char_11,
        input [7:0] char_12,
        input [7:0] char_13,
        input [7:0] char_14,
        input [7:0] char_15,
        input [7:0] char_16,
        input [7:0] char_17,
        input [7:0] char_18,
        input [7:0] char_19,
        input [7:0] char_20,
        input [7:0] char_21,
        input [7:0] char_22,
        input [7:0] char_23,
        input [7:0] char_24,
        input [7:0] char_25,
        input [7:0] char_26,
        input [7:0] char_27,
        input [7:0] char_28,
        input [7:0] char_29,
        input [7:0] char_30,
        input [7:0] char_31,
        input [7:0] char_32,
        input [7:0] char_33,
        input [7:0] char_34,
        input [7:0] char_35,
        input [7:0] char_36,

        input   [9:0]       pixel_x,
        input   [9:0]       pixel_y,
        input               video_on,
        input               vga_clk,

        output  reg     [3:0]       vga_r,
        output  reg     [3:0]       vga_g,
        output  reg     [3:0]       vga_b        
    );


    	// 显示器可显示区域
	// parameter UP_BOUND = 31;
	// parameter DOWN_BOUND = 510;
	parameter LEFT_BOUND = 4;
	parameter RIGHT_BOUND = 783;
    
    parameter left_pos = 144;
    parameter right_pos = 783;

    parameter up_pos_row1 = 31;
    parameter down_pos_row1 = 100;

    parameter up_pos_row2 = 111;
    parameter down_pos_row2 = 180;

    parameter up_pos_row3 = 191;
    parameter down_pos_row3 = 260;

	wire [69:0] row1 [639:0];
    wire [69:0] row2 [639:0];
    wire [69:0] row3 [639:0];

vga_gen_col col_row1_char1(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_1),
	.col_reg_0(row1[5]),
	.col_reg_1(row1[6]),
	.col_reg_2(row1[7]),
	.col_reg_3(row1[8]),
	.col_reg_4(row1[9]),
	.col_reg_5(row1[10]),
	.col_reg_6(row1[11]),
	.col_reg_7(row1[12]),
	.col_reg_8(row1[13]),
	.col_reg_9(row1[14]),
	.col_reg_10(row1[15]),
	.col_reg_11(row1[16]),
	.col_reg_12(row1[17]),
	.col_reg_13(row1[18]),
	.col_reg_14(row1[19]),
	.col_reg_15(row1[20]),
	.col_reg_16(row1[21]),
	.col_reg_17(row1[22]),
	.col_reg_18(row1[23]),
	.col_reg_19(row1[24]),
	.col_reg_20(row1[25]),
	.col_reg_21(row1[26]),
	.col_reg_22(row1[27]),
	.col_reg_23(row1[28]),
	.col_reg_24(row1[29]),
	.col_reg_25(row1[30]),
	.col_reg_26(row1[31]),
	.col_reg_27(row1[32]),
	.col_reg_28(row1[33]),
	.col_reg_29(row1[34]),
	.col_reg_30(row1[35]),
	.col_reg_31(row1[36]),
	.col_reg_32(row1[37]),
	.col_reg_33(row1[38]),
	.col_reg_34(row1[39]),
	.col_reg_35(row1[40]),
	.col_reg_36(row1[41]),
	.col_reg_37(row1[42]),
	.col_reg_38(row1[43]),
	.col_reg_39(row1[44]),
	.col_reg_40(row1[45]),
	.col_reg_41(row1[46]),
	.col_reg_42(row1[47]),
	.col_reg_43(row1[48]),
	.col_reg_44(row1[49]),
	.col_reg_45(row1[50]),
	.col_reg_46(row1[51]),
	.col_reg_47(row1[52]),
	.col_reg_48(row1[53]),
	.col_reg_49(row1[54])
);


vga_gen_col col_row1_char2(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_2),
	.col_reg_0(row1[58]),
	.col_reg_1(row1[59]),
	.col_reg_2(row1[60]),
	.col_reg_3(row1[61]),
	.col_reg_4(row1[62]),
	.col_reg_5(row1[63]),
	.col_reg_6(row1[64]),
	.col_reg_7(row1[65]),
	.col_reg_8(row1[66]),
	.col_reg_9(row1[67]),
	.col_reg_10(row1[68]),
	.col_reg_11(row1[69]),
	.col_reg_12(row1[70]),
	.col_reg_13(row1[71]),
	.col_reg_14(row1[72]),
	.col_reg_15(row1[73]),
	.col_reg_16(row1[74]),
	.col_reg_17(row1[75]),
	.col_reg_18(row1[76]),
	.col_reg_19(row1[77]),
	.col_reg_20(row1[78]),
	.col_reg_21(row1[79]),
	.col_reg_22(row1[80]),
	.col_reg_23(row1[81]),
	.col_reg_24(row1[82]),
	.col_reg_25(row1[83]),
	.col_reg_26(row1[84]),
	.col_reg_27(row1[85]),
	.col_reg_28(row1[86]),
	.col_reg_29(row1[87]),
	.col_reg_30(row1[88]),
	.col_reg_31(row1[89]),
	.col_reg_32(row1[90]),
	.col_reg_33(row1[91]),
	.col_reg_34(row1[92]),
	.col_reg_35(row1[93]),
	.col_reg_36(row1[94]),
	.col_reg_37(row1[95]),
	.col_reg_38(row1[96]),
	.col_reg_39(row1[97]),
	.col_reg_40(row1[98]),
	.col_reg_41(row1[99]),
	.col_reg_42(row1[100]),
	.col_reg_43(row1[101]),
	.col_reg_44(row1[102]),
	.col_reg_45(row1[103]),
	.col_reg_46(row1[104]),
	.col_reg_47(row1[105]),
	.col_reg_48(row1[106]),
	.col_reg_49(row1[107])
);


vga_gen_col col_row1_char3(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_3),
	.col_reg_0(row1[111]),
	.col_reg_1(row1[112]),
	.col_reg_2(row1[113]),
	.col_reg_3(row1[114]),
	.col_reg_4(row1[115]),
	.col_reg_5(row1[116]),
	.col_reg_6(row1[117]),
	.col_reg_7(row1[118]),
	.col_reg_8(row1[119]),
	.col_reg_9(row1[120]),
	.col_reg_10(row1[121]),
	.col_reg_11(row1[122]),
	.col_reg_12(row1[123]),
	.col_reg_13(row1[124]),
	.col_reg_14(row1[125]),
	.col_reg_15(row1[126]),
	.col_reg_16(row1[127]),
	.col_reg_17(row1[128]),
	.col_reg_18(row1[129]),
	.col_reg_19(row1[130]),
	.col_reg_20(row1[131]),
	.col_reg_21(row1[132]),
	.col_reg_22(row1[133]),
	.col_reg_23(row1[134]),
	.col_reg_24(row1[135]),
	.col_reg_25(row1[136]),
	.col_reg_26(row1[137]),
	.col_reg_27(row1[138]),
	.col_reg_28(row1[139]),
	.col_reg_29(row1[140]),
	.col_reg_30(row1[141]),
	.col_reg_31(row1[142]),
	.col_reg_32(row1[143]),
	.col_reg_33(row1[144]),
	.col_reg_34(row1[145]),
	.col_reg_35(row1[146]),
	.col_reg_36(row1[147]),
	.col_reg_37(row1[148]),
	.col_reg_38(row1[149]),
	.col_reg_39(row1[150]),
	.col_reg_40(row1[151]),
	.col_reg_41(row1[152]),
	.col_reg_42(row1[153]),
	.col_reg_43(row1[154]),
	.col_reg_44(row1[155]),
	.col_reg_45(row1[156]),
	.col_reg_46(row1[157]),
	.col_reg_47(row1[158]),
	.col_reg_48(row1[159]),
	.col_reg_49(row1[160])
);


vga_gen_col col_row1_char4(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_4),
	.col_reg_0(row1[164]),
	.col_reg_1(row1[165]),
	.col_reg_2(row1[166]),
	.col_reg_3(row1[167]),
	.col_reg_4(row1[168]),
	.col_reg_5(row1[169]),
	.col_reg_6(row1[170]),
	.col_reg_7(row1[171]),
	.col_reg_8(row1[172]),
	.col_reg_9(row1[173]),
	.col_reg_10(row1[174]),
	.col_reg_11(row1[175]),
	.col_reg_12(row1[176]),
	.col_reg_13(row1[177]),
	.col_reg_14(row1[178]),
	.col_reg_15(row1[179]),
	.col_reg_16(row1[180]),
	.col_reg_17(row1[181]),
	.col_reg_18(row1[182]),
	.col_reg_19(row1[183]),
	.col_reg_20(row1[184]),
	.col_reg_21(row1[185]),
	.col_reg_22(row1[186]),
	.col_reg_23(row1[187]),
	.col_reg_24(row1[188]),
	.col_reg_25(row1[189]),
	.col_reg_26(row1[190]),
	.col_reg_27(row1[191]),
	.col_reg_28(row1[192]),
	.col_reg_29(row1[193]),
	.col_reg_30(row1[194]),
	.col_reg_31(row1[195]),
	.col_reg_32(row1[196]),
	.col_reg_33(row1[197]),
	.col_reg_34(row1[198]),
	.col_reg_35(row1[199]),
	.col_reg_36(row1[200]),
	.col_reg_37(row1[201]),
	.col_reg_38(row1[202]),
	.col_reg_39(row1[203]),
	.col_reg_40(row1[204]),
	.col_reg_41(row1[205]),
	.col_reg_42(row1[206]),
	.col_reg_43(row1[207]),
	.col_reg_44(row1[208]),
	.col_reg_45(row1[209]),
	.col_reg_46(row1[210]),
	.col_reg_47(row1[211]),
	.col_reg_48(row1[212]),
	.col_reg_49(row1[213])
);


vga_gen_col col_row1_char5(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_5),
	.col_reg_0(row1[217]),
	.col_reg_1(row1[218]),
	.col_reg_2(row1[219]),
	.col_reg_3(row1[220]),
	.col_reg_4(row1[221]),
	.col_reg_5(row1[222]),
	.col_reg_6(row1[223]),
	.col_reg_7(row1[224]),
	.col_reg_8(row1[225]),
	.col_reg_9(row1[226]),
	.col_reg_10(row1[227]),
	.col_reg_11(row1[228]),
	.col_reg_12(row1[229]),
	.col_reg_13(row1[230]),
	.col_reg_14(row1[231]),
	.col_reg_15(row1[232]),
	.col_reg_16(row1[233]),
	.col_reg_17(row1[234]),
	.col_reg_18(row1[235]),
	.col_reg_19(row1[236]),
	.col_reg_20(row1[237]),
	.col_reg_21(row1[238]),
	.col_reg_22(row1[239]),
	.col_reg_23(row1[240]),
	.col_reg_24(row1[241]),
	.col_reg_25(row1[242]),
	.col_reg_26(row1[243]),
	.col_reg_27(row1[244]),
	.col_reg_28(row1[245]),
	.col_reg_29(row1[246]),
	.col_reg_30(row1[247]),
	.col_reg_31(row1[248]),
	.col_reg_32(row1[249]),
	.col_reg_33(row1[250]),
	.col_reg_34(row1[251]),
	.col_reg_35(row1[252]),
	.col_reg_36(row1[253]),
	.col_reg_37(row1[254]),
	.col_reg_38(row1[255]),
	.col_reg_39(row1[256]),
	.col_reg_40(row1[257]),
	.col_reg_41(row1[258]),
	.col_reg_42(row1[259]),
	.col_reg_43(row1[260]),
	.col_reg_44(row1[261]),
	.col_reg_45(row1[262]),
	.col_reg_46(row1[263]),
	.col_reg_47(row1[264]),
	.col_reg_48(row1[265]),
	.col_reg_49(row1[266])
);


vga_gen_col col_row1_char6(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_6),
	.col_reg_0(row1[270]),
	.col_reg_1(row1[271]),
	.col_reg_2(row1[272]),
	.col_reg_3(row1[273]),
	.col_reg_4(row1[274]),
	.col_reg_5(row1[275]),
	.col_reg_6(row1[276]),
	.col_reg_7(row1[277]),
	.col_reg_8(row1[278]),
	.col_reg_9(row1[279]),
	.col_reg_10(row1[280]),
	.col_reg_11(row1[281]),
	.col_reg_12(row1[282]),
	.col_reg_13(row1[283]),
	.col_reg_14(row1[284]),
	.col_reg_15(row1[285]),
	.col_reg_16(row1[286]),
	.col_reg_17(row1[287]),
	.col_reg_18(row1[288]),
	.col_reg_19(row1[289]),
	.col_reg_20(row1[290]),
	.col_reg_21(row1[291]),
	.col_reg_22(row1[292]),
	.col_reg_23(row1[293]),
	.col_reg_24(row1[294]),
	.col_reg_25(row1[295]),
	.col_reg_26(row1[296]),
	.col_reg_27(row1[297]),
	.col_reg_28(row1[298]),
	.col_reg_29(row1[299]),
	.col_reg_30(row1[300]),
	.col_reg_31(row1[301]),
	.col_reg_32(row1[302]),
	.col_reg_33(row1[303]),
	.col_reg_34(row1[304]),
	.col_reg_35(row1[305]),
	.col_reg_36(row1[306]),
	.col_reg_37(row1[307]),
	.col_reg_38(row1[308]),
	.col_reg_39(row1[309]),
	.col_reg_40(row1[310]),
	.col_reg_41(row1[311]),
	.col_reg_42(row1[312]),
	.col_reg_43(row1[313]),
	.col_reg_44(row1[314]),
	.col_reg_45(row1[315]),
	.col_reg_46(row1[316]),
	.col_reg_47(row1[317]),
	.col_reg_48(row1[318]),
	.col_reg_49(row1[319])
);


vga_gen_col col_row1_char7(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_7),
	.col_reg_0(row1[323]),
	.col_reg_1(row1[324]),
	.col_reg_2(row1[325]),
	.col_reg_3(row1[326]),
	.col_reg_4(row1[327]),
	.col_reg_5(row1[328]),
	.col_reg_6(row1[329]),
	.col_reg_7(row1[330]),
	.col_reg_8(row1[331]),
	.col_reg_9(row1[332]),
	.col_reg_10(row1[333]),
	.col_reg_11(row1[334]),
	.col_reg_12(row1[335]),
	.col_reg_13(row1[336]),
	.col_reg_14(row1[337]),
	.col_reg_15(row1[338]),
	.col_reg_16(row1[339]),
	.col_reg_17(row1[340]),
	.col_reg_18(row1[341]),
	.col_reg_19(row1[342]),
	.col_reg_20(row1[343]),
	.col_reg_21(row1[344]),
	.col_reg_22(row1[345]),
	.col_reg_23(row1[346]),
	.col_reg_24(row1[347]),
	.col_reg_25(row1[348]),
	.col_reg_26(row1[349]),
	.col_reg_27(row1[350]),
	.col_reg_28(row1[351]),
	.col_reg_29(row1[352]),
	.col_reg_30(row1[353]),
	.col_reg_31(row1[354]),
	.col_reg_32(row1[355]),
	.col_reg_33(row1[356]),
	.col_reg_34(row1[357]),
	.col_reg_35(row1[358]),
	.col_reg_36(row1[359]),
	.col_reg_37(row1[360]),
	.col_reg_38(row1[361]),
	.col_reg_39(row1[362]),
	.col_reg_40(row1[363]),
	.col_reg_41(row1[364]),
	.col_reg_42(row1[365]),
	.col_reg_43(row1[366]),
	.col_reg_44(row1[367]),
	.col_reg_45(row1[368]),
	.col_reg_46(row1[369]),
	.col_reg_47(row1[370]),
	.col_reg_48(row1[371]),
	.col_reg_49(row1[372])
);


vga_gen_col col_row1_char8(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_8),
	.col_reg_0(row1[376]),
	.col_reg_1(row1[377]),
	.col_reg_2(row1[378]),
	.col_reg_3(row1[379]),
	.col_reg_4(row1[380]),
	.col_reg_5(row1[381]),
	.col_reg_6(row1[382]),
	.col_reg_7(row1[383]),
	.col_reg_8(row1[384]),
	.col_reg_9(row1[385]),
	.col_reg_10(row1[386]),
	.col_reg_11(row1[387]),
	.col_reg_12(row1[388]),
	.col_reg_13(row1[389]),
	.col_reg_14(row1[390]),
	.col_reg_15(row1[391]),
	.col_reg_16(row1[392]),
	.col_reg_17(row1[393]),
	.col_reg_18(row1[394]),
	.col_reg_19(row1[395]),
	.col_reg_20(row1[396]),
	.col_reg_21(row1[397]),
	.col_reg_22(row1[398]),
	.col_reg_23(row1[399]),
	.col_reg_24(row1[400]),
	.col_reg_25(row1[401]),
	.col_reg_26(row1[402]),
	.col_reg_27(row1[403]),
	.col_reg_28(row1[404]),
	.col_reg_29(row1[405]),
	.col_reg_30(row1[406]),
	.col_reg_31(row1[407]),
	.col_reg_32(row1[408]),
	.col_reg_33(row1[409]),
	.col_reg_34(row1[410]),
	.col_reg_35(row1[411]),
	.col_reg_36(row1[412]),
	.col_reg_37(row1[413]),
	.col_reg_38(row1[414]),
	.col_reg_39(row1[415]),
	.col_reg_40(row1[416]),
	.col_reg_41(row1[417]),
	.col_reg_42(row1[418]),
	.col_reg_43(row1[419]),
	.col_reg_44(row1[420]),
	.col_reg_45(row1[421]),
	.col_reg_46(row1[422]),
	.col_reg_47(row1[423]),
	.col_reg_48(row1[424]),
	.col_reg_49(row1[425])
);


vga_gen_col col_row1_char9(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_9),
	.col_reg_0(row1[429]),
	.col_reg_1(row1[430]),
	.col_reg_2(row1[431]),
	.col_reg_3(row1[432]),
	.col_reg_4(row1[433]),
	.col_reg_5(row1[434]),
	.col_reg_6(row1[435]),
	.col_reg_7(row1[436]),
	.col_reg_8(row1[437]),
	.col_reg_9(row1[438]),
	.col_reg_10(row1[439]),
	.col_reg_11(row1[440]),
	.col_reg_12(row1[441]),
	.col_reg_13(row1[442]),
	.col_reg_14(row1[443]),
	.col_reg_15(row1[444]),
	.col_reg_16(row1[445]),
	.col_reg_17(row1[446]),
	.col_reg_18(row1[447]),
	.col_reg_19(row1[448]),
	.col_reg_20(row1[449]),
	.col_reg_21(row1[450]),
	.col_reg_22(row1[451]),
	.col_reg_23(row1[452]),
	.col_reg_24(row1[453]),
	.col_reg_25(row1[454]),
	.col_reg_26(row1[455]),
	.col_reg_27(row1[456]),
	.col_reg_28(row1[457]),
	.col_reg_29(row1[458]),
	.col_reg_30(row1[459]),
	.col_reg_31(row1[460]),
	.col_reg_32(row1[461]),
	.col_reg_33(row1[462]),
	.col_reg_34(row1[463]),
	.col_reg_35(row1[464]),
	.col_reg_36(row1[465]),
	.col_reg_37(row1[466]),
	.col_reg_38(row1[467]),
	.col_reg_39(row1[468]),
	.col_reg_40(row1[469]),
	.col_reg_41(row1[470]),
	.col_reg_42(row1[471]),
	.col_reg_43(row1[472]),
	.col_reg_44(row1[473]),
	.col_reg_45(row1[474]),
	.col_reg_46(row1[475]),
	.col_reg_47(row1[476]),
	.col_reg_48(row1[477]),
	.col_reg_49(row1[478])
);


vga_gen_col col_row1_char10(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_10),
	.col_reg_0(row1[482]),
	.col_reg_1(row1[483]),
	.col_reg_2(row1[484]),
	.col_reg_3(row1[485]),
	.col_reg_4(row1[486]),
	.col_reg_5(row1[487]),
	.col_reg_6(row1[488]),
	.col_reg_7(row1[489]),
	.col_reg_8(row1[490]),
	.col_reg_9(row1[491]),
	.col_reg_10(row1[492]),
	.col_reg_11(row1[493]),
	.col_reg_12(row1[494]),
	.col_reg_13(row1[495]),
	.col_reg_14(row1[496]),
	.col_reg_15(row1[497]),
	.col_reg_16(row1[498]),
	.col_reg_17(row1[499]),
	.col_reg_18(row1[500]),
	.col_reg_19(row1[501]),
	.col_reg_20(row1[502]),
	.col_reg_21(row1[503]),
	.col_reg_22(row1[504]),
	.col_reg_23(row1[505]),
	.col_reg_24(row1[506]),
	.col_reg_25(row1[507]),
	.col_reg_26(row1[508]),
	.col_reg_27(row1[509]),
	.col_reg_28(row1[510]),
	.col_reg_29(row1[511]),
	.col_reg_30(row1[512]),
	.col_reg_31(row1[513]),
	.col_reg_32(row1[514]),
	.col_reg_33(row1[515]),
	.col_reg_34(row1[516]),
	.col_reg_35(row1[517]),
	.col_reg_36(row1[518]),
	.col_reg_37(row1[519]),
	.col_reg_38(row1[520]),
	.col_reg_39(row1[521]),
	.col_reg_40(row1[522]),
	.col_reg_41(row1[523]),
	.col_reg_42(row1[524]),
	.col_reg_43(row1[525]),
	.col_reg_44(row1[526]),
	.col_reg_45(row1[527]),
	.col_reg_46(row1[528]),
	.col_reg_47(row1[529]),
	.col_reg_48(row1[530]),
	.col_reg_49(row1[531])
);


vga_gen_col col_row1_char11(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_11),
	.col_reg_0(row1[535]),
	.col_reg_1(row1[536]),
	.col_reg_2(row1[537]),
	.col_reg_3(row1[538]),
	.col_reg_4(row1[539]),
	.col_reg_5(row1[540]),
	.col_reg_6(row1[541]),
	.col_reg_7(row1[542]),
	.col_reg_8(row1[543]),
	.col_reg_9(row1[544]),
	.col_reg_10(row1[545]),
	.col_reg_11(row1[546]),
	.col_reg_12(row1[547]),
	.col_reg_13(row1[548]),
	.col_reg_14(row1[549]),
	.col_reg_15(row1[550]),
	.col_reg_16(row1[551]),
	.col_reg_17(row1[552]),
	.col_reg_18(row1[553]),
	.col_reg_19(row1[554]),
	.col_reg_20(row1[555]),
	.col_reg_21(row1[556]),
	.col_reg_22(row1[557]),
	.col_reg_23(row1[558]),
	.col_reg_24(row1[559]),
	.col_reg_25(row1[560]),
	.col_reg_26(row1[561]),
	.col_reg_27(row1[562]),
	.col_reg_28(row1[563]),
	.col_reg_29(row1[564]),
	.col_reg_30(row1[565]),
	.col_reg_31(row1[566]),
	.col_reg_32(row1[567]),
	.col_reg_33(row1[568]),
	.col_reg_34(row1[569]),
	.col_reg_35(row1[570]),
	.col_reg_36(row1[571]),
	.col_reg_37(row1[572]),
	.col_reg_38(row1[573]),
	.col_reg_39(row1[574]),
	.col_reg_40(row1[575]),
	.col_reg_41(row1[576]),
	.col_reg_42(row1[577]),
	.col_reg_43(row1[578]),
	.col_reg_44(row1[579]),
	.col_reg_45(row1[580]),
	.col_reg_46(row1[581]),
	.col_reg_47(row1[582]),
	.col_reg_48(row1[583]),
	.col_reg_49(row1[584])
);


vga_gen_col col_row1_char12(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_12),
	.col_reg_0(row1[588]),
	.col_reg_1(row1[589]),
	.col_reg_2(row1[590]),
	.col_reg_3(row1[591]),
	.col_reg_4(row1[592]),
	.col_reg_5(row1[593]),
	.col_reg_6(row1[594]),
	.col_reg_7(row1[595]),
	.col_reg_8(row1[596]),
	.col_reg_9(row1[597]),
	.col_reg_10(row1[598]),
	.col_reg_11(row1[599]),
	.col_reg_12(row1[600]),
	.col_reg_13(row1[601]),
	.col_reg_14(row1[602]),
	.col_reg_15(row1[603]),
	.col_reg_16(row1[604]),
	.col_reg_17(row1[605]),
	.col_reg_18(row1[606]),
	.col_reg_19(row1[607]),
	.col_reg_20(row1[608]),
	.col_reg_21(row1[609]),
	.col_reg_22(row1[610]),
	.col_reg_23(row1[611]),
	.col_reg_24(row1[612]),
	.col_reg_25(row1[613]),
	.col_reg_26(row1[614]),
	.col_reg_27(row1[615]),
	.col_reg_28(row1[616]),
	.col_reg_29(row1[617]),
	.col_reg_30(row1[618]),
	.col_reg_31(row1[619]),
	.col_reg_32(row1[620]),
	.col_reg_33(row1[621]),
	.col_reg_34(row1[622]),
	.col_reg_35(row1[623]),
	.col_reg_36(row1[624]),
	.col_reg_37(row1[625]),
	.col_reg_38(row1[626]),
	.col_reg_39(row1[627]),
	.col_reg_40(row1[628]),
	.col_reg_41(row1[629]),
	.col_reg_42(row1[630]),
	.col_reg_43(row1[631]),
	.col_reg_44(row1[632]),
	.col_reg_45(row1[633]),
	.col_reg_46(row1[634]),
	.col_reg_47(row1[635]),
	.col_reg_48(row1[636]),
	.col_reg_49(row1[637])
);


vga_gen_col col_row2_char1(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_13),
	.col_reg_0(row2[5]),
	.col_reg_1(row2[6]),
	.col_reg_2(row2[7]),
	.col_reg_3(row2[8]),
	.col_reg_4(row2[9]),
	.col_reg_5(row2[10]),
	.col_reg_6(row2[11]),
	.col_reg_7(row2[12]),
	.col_reg_8(row2[13]),
	.col_reg_9(row2[14]),
	.col_reg_10(row2[15]),
	.col_reg_11(row2[16]),
	.col_reg_12(row2[17]),
	.col_reg_13(row2[18]),
	.col_reg_14(row2[19]),
	.col_reg_15(row2[20]),
	.col_reg_16(row2[21]),
	.col_reg_17(row2[22]),
	.col_reg_18(row2[23]),
	.col_reg_19(row2[24]),
	.col_reg_20(row2[25]),
	.col_reg_21(row2[26]),
	.col_reg_22(row2[27]),
	.col_reg_23(row2[28]),
	.col_reg_24(row2[29]),
	.col_reg_25(row2[30]),
	.col_reg_26(row2[31]),
	.col_reg_27(row2[32]),
	.col_reg_28(row2[33]),
	.col_reg_29(row2[34]),
	.col_reg_30(row2[35]),
	.col_reg_31(row2[36]),
	.col_reg_32(row2[37]),
	.col_reg_33(row2[38]),
	.col_reg_34(row2[39]),
	.col_reg_35(row2[40]),
	.col_reg_36(row2[41]),
	.col_reg_37(row2[42]),
	.col_reg_38(row2[43]),
	.col_reg_39(row2[44]),
	.col_reg_40(row2[45]),
	.col_reg_41(row2[46]),
	.col_reg_42(row2[47]),
	.col_reg_43(row2[48]),
	.col_reg_44(row2[49]),
	.col_reg_45(row2[50]),
	.col_reg_46(row2[51]),
	.col_reg_47(row2[52]),
	.col_reg_48(row2[53]),
	.col_reg_49(row2[54])
);


vga_gen_col col_row2_char2(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_14),
	.col_reg_0(row2[58]),
	.col_reg_1(row2[59]),
	.col_reg_2(row2[60]),
	.col_reg_3(row2[61]),
	.col_reg_4(row2[62]),
	.col_reg_5(row2[63]),
	.col_reg_6(row2[64]),
	.col_reg_7(row2[65]),
	.col_reg_8(row2[66]),
	.col_reg_9(row2[67]),
	.col_reg_10(row2[68]),
	.col_reg_11(row2[69]),
	.col_reg_12(row2[70]),
	.col_reg_13(row2[71]),
	.col_reg_14(row2[72]),
	.col_reg_15(row2[73]),
	.col_reg_16(row2[74]),
	.col_reg_17(row2[75]),
	.col_reg_18(row2[76]),
	.col_reg_19(row2[77]),
	.col_reg_20(row2[78]),
	.col_reg_21(row2[79]),
	.col_reg_22(row2[80]),
	.col_reg_23(row2[81]),
	.col_reg_24(row2[82]),
	.col_reg_25(row2[83]),
	.col_reg_26(row2[84]),
	.col_reg_27(row2[85]),
	.col_reg_28(row2[86]),
	.col_reg_29(row2[87]),
	.col_reg_30(row2[88]),
	.col_reg_31(row2[89]),
	.col_reg_32(row2[90]),
	.col_reg_33(row2[91]),
	.col_reg_34(row2[92]),
	.col_reg_35(row2[93]),
	.col_reg_36(row2[94]),
	.col_reg_37(row2[95]),
	.col_reg_38(row2[96]),
	.col_reg_39(row2[97]),
	.col_reg_40(row2[98]),
	.col_reg_41(row2[99]),
	.col_reg_42(row2[100]),
	.col_reg_43(row2[101]),
	.col_reg_44(row2[102]),
	.col_reg_45(row2[103]),
	.col_reg_46(row2[104]),
	.col_reg_47(row2[105]),
	.col_reg_48(row2[106]),
	.col_reg_49(row2[107])
);


vga_gen_col col_row2_char3(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_15),
	.col_reg_0(row2[111]),
	.col_reg_1(row2[112]),
	.col_reg_2(row2[113]),
	.col_reg_3(row2[114]),
	.col_reg_4(row2[115]),
	.col_reg_5(row2[116]),
	.col_reg_6(row2[117]),
	.col_reg_7(row2[118]),
	.col_reg_8(row2[119]),
	.col_reg_9(row2[120]),
	.col_reg_10(row2[121]),
	.col_reg_11(row2[122]),
	.col_reg_12(row2[123]),
	.col_reg_13(row2[124]),
	.col_reg_14(row2[125]),
	.col_reg_15(row2[126]),
	.col_reg_16(row2[127]),
	.col_reg_17(row2[128]),
	.col_reg_18(row2[129]),
	.col_reg_19(row2[130]),
	.col_reg_20(row2[131]),
	.col_reg_21(row2[132]),
	.col_reg_22(row2[133]),
	.col_reg_23(row2[134]),
	.col_reg_24(row2[135]),
	.col_reg_25(row2[136]),
	.col_reg_26(row2[137]),
	.col_reg_27(row2[138]),
	.col_reg_28(row2[139]),
	.col_reg_29(row2[140]),
	.col_reg_30(row2[141]),
	.col_reg_31(row2[142]),
	.col_reg_32(row2[143]),
	.col_reg_33(row2[144]),
	.col_reg_34(row2[145]),
	.col_reg_35(row2[146]),
	.col_reg_36(row2[147]),
	.col_reg_37(row2[148]),
	.col_reg_38(row2[149]),
	.col_reg_39(row2[150]),
	.col_reg_40(row2[151]),
	.col_reg_41(row2[152]),
	.col_reg_42(row2[153]),
	.col_reg_43(row2[154]),
	.col_reg_44(row2[155]),
	.col_reg_45(row2[156]),
	.col_reg_46(row2[157]),
	.col_reg_47(row2[158]),
	.col_reg_48(row2[159]),
	.col_reg_49(row2[160])
);


vga_gen_col col_row2_char4(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_16),
	.col_reg_0(row2[164]),
	.col_reg_1(row2[165]),
	.col_reg_2(row2[166]),
	.col_reg_3(row2[167]),
	.col_reg_4(row2[168]),
	.col_reg_5(row2[169]),
	.col_reg_6(row2[170]),
	.col_reg_7(row2[171]),
	.col_reg_8(row2[172]),
	.col_reg_9(row2[173]),
	.col_reg_10(row2[174]),
	.col_reg_11(row2[175]),
	.col_reg_12(row2[176]),
	.col_reg_13(row2[177]),
	.col_reg_14(row2[178]),
	.col_reg_15(row2[179]),
	.col_reg_16(row2[180]),
	.col_reg_17(row2[181]),
	.col_reg_18(row2[182]),
	.col_reg_19(row2[183]),
	.col_reg_20(row2[184]),
	.col_reg_21(row2[185]),
	.col_reg_22(row2[186]),
	.col_reg_23(row2[187]),
	.col_reg_24(row2[188]),
	.col_reg_25(row2[189]),
	.col_reg_26(row2[190]),
	.col_reg_27(row2[191]),
	.col_reg_28(row2[192]),
	.col_reg_29(row2[193]),
	.col_reg_30(row2[194]),
	.col_reg_31(row2[195]),
	.col_reg_32(row2[196]),
	.col_reg_33(row2[197]),
	.col_reg_34(row2[198]),
	.col_reg_35(row2[199]),
	.col_reg_36(row2[200]),
	.col_reg_37(row2[201]),
	.col_reg_38(row2[202]),
	.col_reg_39(row2[203]),
	.col_reg_40(row2[204]),
	.col_reg_41(row2[205]),
	.col_reg_42(row2[206]),
	.col_reg_43(row2[207]),
	.col_reg_44(row2[208]),
	.col_reg_45(row2[209]),
	.col_reg_46(row2[210]),
	.col_reg_47(row2[211]),
	.col_reg_48(row2[212]),
	.col_reg_49(row2[213])
);


vga_gen_col col_row2_char5(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_17),
	.col_reg_0(row2[217]),
	.col_reg_1(row2[218]),
	.col_reg_2(row2[219]),
	.col_reg_3(row2[220]),
	.col_reg_4(row2[221]),
	.col_reg_5(row2[222]),
	.col_reg_6(row2[223]),
	.col_reg_7(row2[224]),
	.col_reg_8(row2[225]),
	.col_reg_9(row2[226]),
	.col_reg_10(row2[227]),
	.col_reg_11(row2[228]),
	.col_reg_12(row2[229]),
	.col_reg_13(row2[230]),
	.col_reg_14(row2[231]),
	.col_reg_15(row2[232]),
	.col_reg_16(row2[233]),
	.col_reg_17(row2[234]),
	.col_reg_18(row2[235]),
	.col_reg_19(row2[236]),
	.col_reg_20(row2[237]),
	.col_reg_21(row2[238]),
	.col_reg_22(row2[239]),
	.col_reg_23(row2[240]),
	.col_reg_24(row2[241]),
	.col_reg_25(row2[242]),
	.col_reg_26(row2[243]),
	.col_reg_27(row2[244]),
	.col_reg_28(row2[245]),
	.col_reg_29(row2[246]),
	.col_reg_30(row2[247]),
	.col_reg_31(row2[248]),
	.col_reg_32(row2[249]),
	.col_reg_33(row2[250]),
	.col_reg_34(row2[251]),
	.col_reg_35(row2[252]),
	.col_reg_36(row2[253]),
	.col_reg_37(row2[254]),
	.col_reg_38(row2[255]),
	.col_reg_39(row2[256]),
	.col_reg_40(row2[257]),
	.col_reg_41(row2[258]),
	.col_reg_42(row2[259]),
	.col_reg_43(row2[260]),
	.col_reg_44(row2[261]),
	.col_reg_45(row2[262]),
	.col_reg_46(row2[263]),
	.col_reg_47(row2[264]),
	.col_reg_48(row2[265]),
	.col_reg_49(row2[266])
);


vga_gen_col col_row2_char6(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_18),
	.col_reg_0(row2[270]),
	.col_reg_1(row2[271]),
	.col_reg_2(row2[272]),
	.col_reg_3(row2[273]),
	.col_reg_4(row2[274]),
	.col_reg_5(row2[275]),
	.col_reg_6(row2[276]),
	.col_reg_7(row2[277]),
	.col_reg_8(row2[278]),
	.col_reg_9(row2[279]),
	.col_reg_10(row2[280]),
	.col_reg_11(row2[281]),
	.col_reg_12(row2[282]),
	.col_reg_13(row2[283]),
	.col_reg_14(row2[284]),
	.col_reg_15(row2[285]),
	.col_reg_16(row2[286]),
	.col_reg_17(row2[287]),
	.col_reg_18(row2[288]),
	.col_reg_19(row2[289]),
	.col_reg_20(row2[290]),
	.col_reg_21(row2[291]),
	.col_reg_22(row2[292]),
	.col_reg_23(row2[293]),
	.col_reg_24(row2[294]),
	.col_reg_25(row2[295]),
	.col_reg_26(row2[296]),
	.col_reg_27(row2[297]),
	.col_reg_28(row2[298]),
	.col_reg_29(row2[299]),
	.col_reg_30(row2[300]),
	.col_reg_31(row2[301]),
	.col_reg_32(row2[302]),
	.col_reg_33(row2[303]),
	.col_reg_34(row2[304]),
	.col_reg_35(row2[305]),
	.col_reg_36(row2[306]),
	.col_reg_37(row2[307]),
	.col_reg_38(row2[308]),
	.col_reg_39(row2[309]),
	.col_reg_40(row2[310]),
	.col_reg_41(row2[311]),
	.col_reg_42(row2[312]),
	.col_reg_43(row2[313]),
	.col_reg_44(row2[314]),
	.col_reg_45(row2[315]),
	.col_reg_46(row2[316]),
	.col_reg_47(row2[317]),
	.col_reg_48(row2[318]),
	.col_reg_49(row2[319])
);


vga_gen_col col_row2_char7(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_19),
	.col_reg_0(row2[323]),
	.col_reg_1(row2[324]),
	.col_reg_2(row2[325]),
	.col_reg_3(row2[326]),
	.col_reg_4(row2[327]),
	.col_reg_5(row2[328]),
	.col_reg_6(row2[329]),
	.col_reg_7(row2[330]),
	.col_reg_8(row2[331]),
	.col_reg_9(row2[332]),
	.col_reg_10(row2[333]),
	.col_reg_11(row2[334]),
	.col_reg_12(row2[335]),
	.col_reg_13(row2[336]),
	.col_reg_14(row2[337]),
	.col_reg_15(row2[338]),
	.col_reg_16(row2[339]),
	.col_reg_17(row2[340]),
	.col_reg_18(row2[341]),
	.col_reg_19(row2[342]),
	.col_reg_20(row2[343]),
	.col_reg_21(row2[344]),
	.col_reg_22(row2[345]),
	.col_reg_23(row2[346]),
	.col_reg_24(row2[347]),
	.col_reg_25(row2[348]),
	.col_reg_26(row2[349]),
	.col_reg_27(row2[350]),
	.col_reg_28(row2[351]),
	.col_reg_29(row2[352]),
	.col_reg_30(row2[353]),
	.col_reg_31(row2[354]),
	.col_reg_32(row2[355]),
	.col_reg_33(row2[356]),
	.col_reg_34(row2[357]),
	.col_reg_35(row2[358]),
	.col_reg_36(row2[359]),
	.col_reg_37(row2[360]),
	.col_reg_38(row2[361]),
	.col_reg_39(row2[362]),
	.col_reg_40(row2[363]),
	.col_reg_41(row2[364]),
	.col_reg_42(row2[365]),
	.col_reg_43(row2[366]),
	.col_reg_44(row2[367]),
	.col_reg_45(row2[368]),
	.col_reg_46(row2[369]),
	.col_reg_47(row2[370]),
	.col_reg_48(row2[371]),
	.col_reg_49(row2[372])
);


vga_gen_col col_row2_char8(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_20),
	.col_reg_0(row2[376]),
	.col_reg_1(row2[377]),
	.col_reg_2(row2[378]),
	.col_reg_3(row2[379]),
	.col_reg_4(row2[380]),
	.col_reg_5(row2[381]),
	.col_reg_6(row2[382]),
	.col_reg_7(row2[383]),
	.col_reg_8(row2[384]),
	.col_reg_9(row2[385]),
	.col_reg_10(row2[386]),
	.col_reg_11(row2[387]),
	.col_reg_12(row2[388]),
	.col_reg_13(row2[389]),
	.col_reg_14(row2[390]),
	.col_reg_15(row2[391]),
	.col_reg_16(row2[392]),
	.col_reg_17(row2[393]),
	.col_reg_18(row2[394]),
	.col_reg_19(row2[395]),
	.col_reg_20(row2[396]),
	.col_reg_21(row2[397]),
	.col_reg_22(row2[398]),
	.col_reg_23(row2[399]),
	.col_reg_24(row2[400]),
	.col_reg_25(row2[401]),
	.col_reg_26(row2[402]),
	.col_reg_27(row2[403]),
	.col_reg_28(row2[404]),
	.col_reg_29(row2[405]),
	.col_reg_30(row2[406]),
	.col_reg_31(row2[407]),
	.col_reg_32(row2[408]),
	.col_reg_33(row2[409]),
	.col_reg_34(row2[410]),
	.col_reg_35(row2[411]),
	.col_reg_36(row2[412]),
	.col_reg_37(row2[413]),
	.col_reg_38(row2[414]),
	.col_reg_39(row2[415]),
	.col_reg_40(row2[416]),
	.col_reg_41(row2[417]),
	.col_reg_42(row2[418]),
	.col_reg_43(row2[419]),
	.col_reg_44(row2[420]),
	.col_reg_45(row2[421]),
	.col_reg_46(row2[422]),
	.col_reg_47(row2[423]),
	.col_reg_48(row2[424]),
	.col_reg_49(row2[425])
);


vga_gen_col col_row2_char9(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_21),
	.col_reg_0(row2[429]),
	.col_reg_1(row2[430]),
	.col_reg_2(row2[431]),
	.col_reg_3(row2[432]),
	.col_reg_4(row2[433]),
	.col_reg_5(row2[434]),
	.col_reg_6(row2[435]),
	.col_reg_7(row2[436]),
	.col_reg_8(row2[437]),
	.col_reg_9(row2[438]),
	.col_reg_10(row2[439]),
	.col_reg_11(row2[440]),
	.col_reg_12(row2[441]),
	.col_reg_13(row2[442]),
	.col_reg_14(row2[443]),
	.col_reg_15(row2[444]),
	.col_reg_16(row2[445]),
	.col_reg_17(row2[446]),
	.col_reg_18(row2[447]),
	.col_reg_19(row2[448]),
	.col_reg_20(row2[449]),
	.col_reg_21(row2[450]),
	.col_reg_22(row2[451]),
	.col_reg_23(row2[452]),
	.col_reg_24(row2[453]),
	.col_reg_25(row2[454]),
	.col_reg_26(row2[455]),
	.col_reg_27(row2[456]),
	.col_reg_28(row2[457]),
	.col_reg_29(row2[458]),
	.col_reg_30(row2[459]),
	.col_reg_31(row2[460]),
	.col_reg_32(row2[461]),
	.col_reg_33(row2[462]),
	.col_reg_34(row2[463]),
	.col_reg_35(row2[464]),
	.col_reg_36(row2[465]),
	.col_reg_37(row2[466]),
	.col_reg_38(row2[467]),
	.col_reg_39(row2[468]),
	.col_reg_40(row2[469]),
	.col_reg_41(row2[470]),
	.col_reg_42(row2[471]),
	.col_reg_43(row2[472]),
	.col_reg_44(row2[473]),
	.col_reg_45(row2[474]),
	.col_reg_46(row2[475]),
	.col_reg_47(row2[476]),
	.col_reg_48(row2[477]),
	.col_reg_49(row2[478])
);


vga_gen_col col_row2_char10(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_22),
	.col_reg_0(row2[482]),
	.col_reg_1(row2[483]),
	.col_reg_2(row2[484]),
	.col_reg_3(row2[485]),
	.col_reg_4(row2[486]),
	.col_reg_5(row2[487]),
	.col_reg_6(row2[488]),
	.col_reg_7(row2[489]),
	.col_reg_8(row2[490]),
	.col_reg_9(row2[491]),
	.col_reg_10(row2[492]),
	.col_reg_11(row2[493]),
	.col_reg_12(row2[494]),
	.col_reg_13(row2[495]),
	.col_reg_14(row2[496]),
	.col_reg_15(row2[497]),
	.col_reg_16(row2[498]),
	.col_reg_17(row2[499]),
	.col_reg_18(row2[500]),
	.col_reg_19(row2[501]),
	.col_reg_20(row2[502]),
	.col_reg_21(row2[503]),
	.col_reg_22(row2[504]),
	.col_reg_23(row2[505]),
	.col_reg_24(row2[506]),
	.col_reg_25(row2[507]),
	.col_reg_26(row2[508]),
	.col_reg_27(row2[509]),
	.col_reg_28(row2[510]),
	.col_reg_29(row2[511]),
	.col_reg_30(row2[512]),
	.col_reg_31(row2[513]),
	.col_reg_32(row2[514]),
	.col_reg_33(row2[515]),
	.col_reg_34(row2[516]),
	.col_reg_35(row2[517]),
	.col_reg_36(row2[518]),
	.col_reg_37(row2[519]),
	.col_reg_38(row2[520]),
	.col_reg_39(row2[521]),
	.col_reg_40(row2[522]),
	.col_reg_41(row2[523]),
	.col_reg_42(row2[524]),
	.col_reg_43(row2[525]),
	.col_reg_44(row2[526]),
	.col_reg_45(row2[527]),
	.col_reg_46(row2[528]),
	.col_reg_47(row2[529]),
	.col_reg_48(row2[530]),
	.col_reg_49(row2[531])
);


vga_gen_col col_row2_char11(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_23),
	.col_reg_0(row2[535]),
	.col_reg_1(row2[536]),
	.col_reg_2(row2[537]),
	.col_reg_3(row2[538]),
	.col_reg_4(row2[539]),
	.col_reg_5(row2[540]),
	.col_reg_6(row2[541]),
	.col_reg_7(row2[542]),
	.col_reg_8(row2[543]),
	.col_reg_9(row2[544]),
	.col_reg_10(row2[545]),
	.col_reg_11(row2[546]),
	.col_reg_12(row2[547]),
	.col_reg_13(row2[548]),
	.col_reg_14(row2[549]),
	.col_reg_15(row2[550]),
	.col_reg_16(row2[551]),
	.col_reg_17(row2[552]),
	.col_reg_18(row2[553]),
	.col_reg_19(row2[554]),
	.col_reg_20(row2[555]),
	.col_reg_21(row2[556]),
	.col_reg_22(row2[557]),
	.col_reg_23(row2[558]),
	.col_reg_24(row2[559]),
	.col_reg_25(row2[560]),
	.col_reg_26(row2[561]),
	.col_reg_27(row2[562]),
	.col_reg_28(row2[563]),
	.col_reg_29(row2[564]),
	.col_reg_30(row2[565]),
	.col_reg_31(row2[566]),
	.col_reg_32(row2[567]),
	.col_reg_33(row2[568]),
	.col_reg_34(row2[569]),
	.col_reg_35(row2[570]),
	.col_reg_36(row2[571]),
	.col_reg_37(row2[572]),
	.col_reg_38(row2[573]),
	.col_reg_39(row2[574]),
	.col_reg_40(row2[575]),
	.col_reg_41(row2[576]),
	.col_reg_42(row2[577]),
	.col_reg_43(row2[578]),
	.col_reg_44(row2[579]),
	.col_reg_45(row2[580]),
	.col_reg_46(row2[581]),
	.col_reg_47(row2[582]),
	.col_reg_48(row2[583]),
	.col_reg_49(row2[584])
);


vga_gen_col col_row2_char12(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_24),
	.col_reg_0(row2[588]),
	.col_reg_1(row2[589]),
	.col_reg_2(row2[590]),
	.col_reg_3(row2[591]),
	.col_reg_4(row2[592]),
	.col_reg_5(row2[593]),
	.col_reg_6(row2[594]),
	.col_reg_7(row2[595]),
	.col_reg_8(row2[596]),
	.col_reg_9(row2[597]),
	.col_reg_10(row2[598]),
	.col_reg_11(row2[599]),
	.col_reg_12(row2[600]),
	.col_reg_13(row2[601]),
	.col_reg_14(row2[602]),
	.col_reg_15(row2[603]),
	.col_reg_16(row2[604]),
	.col_reg_17(row2[605]),
	.col_reg_18(row2[606]),
	.col_reg_19(row2[607]),
	.col_reg_20(row2[608]),
	.col_reg_21(row2[609]),
	.col_reg_22(row2[610]),
	.col_reg_23(row2[611]),
	.col_reg_24(row2[612]),
	.col_reg_25(row2[613]),
	.col_reg_26(row2[614]),
	.col_reg_27(row2[615]),
	.col_reg_28(row2[616]),
	.col_reg_29(row2[617]),
	.col_reg_30(row2[618]),
	.col_reg_31(row2[619]),
	.col_reg_32(row2[620]),
	.col_reg_33(row2[621]),
	.col_reg_34(row2[622]),
	.col_reg_35(row2[623]),
	.col_reg_36(row2[624]),
	.col_reg_37(row2[625]),
	.col_reg_38(row2[626]),
	.col_reg_39(row2[627]),
	.col_reg_40(row2[628]),
	.col_reg_41(row2[629]),
	.col_reg_42(row2[630]),
	.col_reg_43(row2[631]),
	.col_reg_44(row2[632]),
	.col_reg_45(row2[633]),
	.col_reg_46(row2[634]),
	.col_reg_47(row2[635]),
	.col_reg_48(row2[636]),
	.col_reg_49(row2[637])
);


vga_gen_col col_row3_char1(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_25),
	.col_reg_0(row3[5]),
	.col_reg_1(row3[6]),
	.col_reg_2(row3[7]),
	.col_reg_3(row3[8]),
	.col_reg_4(row3[9]),
	.col_reg_5(row3[10]),
	.col_reg_6(row3[11]),
	.col_reg_7(row3[12]),
	.col_reg_8(row3[13]),
	.col_reg_9(row3[14]),
	.col_reg_10(row3[15]),
	.col_reg_11(row3[16]),
	.col_reg_12(row3[17]),
	.col_reg_13(row3[18]),
	.col_reg_14(row3[19]),
	.col_reg_15(row3[20]),
	.col_reg_16(row3[21]),
	.col_reg_17(row3[22]),
	.col_reg_18(row3[23]),
	.col_reg_19(row3[24]),
	.col_reg_20(row3[25]),
	.col_reg_21(row3[26]),
	.col_reg_22(row3[27]),
	.col_reg_23(row3[28]),
	.col_reg_24(row3[29]),
	.col_reg_25(row3[30]),
	.col_reg_26(row3[31]),
	.col_reg_27(row3[32]),
	.col_reg_28(row3[33]),
	.col_reg_29(row3[34]),
	.col_reg_30(row3[35]),
	.col_reg_31(row3[36]),
	.col_reg_32(row3[37]),
	.col_reg_33(row3[38]),
	.col_reg_34(row3[39]),
	.col_reg_35(row3[40]),
	.col_reg_36(row3[41]),
	.col_reg_37(row3[42]),
	.col_reg_38(row3[43]),
	.col_reg_39(row3[44]),
	.col_reg_40(row3[45]),
	.col_reg_41(row3[46]),
	.col_reg_42(row3[47]),
	.col_reg_43(row3[48]),
	.col_reg_44(row3[49]),
	.col_reg_45(row3[50]),
	.col_reg_46(row3[51]),
	.col_reg_47(row3[52]),
	.col_reg_48(row3[53]),
	.col_reg_49(row3[54])
);


vga_gen_col col_row3_char2(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_26),
	.col_reg_0(row3[58]),
	.col_reg_1(row3[59]),
	.col_reg_2(row3[60]),
	.col_reg_3(row3[61]),
	.col_reg_4(row3[62]),
	.col_reg_5(row3[63]),
	.col_reg_6(row3[64]),
	.col_reg_7(row3[65]),
	.col_reg_8(row3[66]),
	.col_reg_9(row3[67]),
	.col_reg_10(row3[68]),
	.col_reg_11(row3[69]),
	.col_reg_12(row3[70]),
	.col_reg_13(row3[71]),
	.col_reg_14(row3[72]),
	.col_reg_15(row3[73]),
	.col_reg_16(row3[74]),
	.col_reg_17(row3[75]),
	.col_reg_18(row3[76]),
	.col_reg_19(row3[77]),
	.col_reg_20(row3[78]),
	.col_reg_21(row3[79]),
	.col_reg_22(row3[80]),
	.col_reg_23(row3[81]),
	.col_reg_24(row3[82]),
	.col_reg_25(row3[83]),
	.col_reg_26(row3[84]),
	.col_reg_27(row3[85]),
	.col_reg_28(row3[86]),
	.col_reg_29(row3[87]),
	.col_reg_30(row3[88]),
	.col_reg_31(row3[89]),
	.col_reg_32(row3[90]),
	.col_reg_33(row3[91]),
	.col_reg_34(row3[92]),
	.col_reg_35(row3[93]),
	.col_reg_36(row3[94]),
	.col_reg_37(row3[95]),
	.col_reg_38(row3[96]),
	.col_reg_39(row3[97]),
	.col_reg_40(row3[98]),
	.col_reg_41(row3[99]),
	.col_reg_42(row3[100]),
	.col_reg_43(row3[101]),
	.col_reg_44(row3[102]),
	.col_reg_45(row3[103]),
	.col_reg_46(row3[104]),
	.col_reg_47(row3[105]),
	.col_reg_48(row3[106]),
	.col_reg_49(row3[107])
);


vga_gen_col col_row3_char3(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_27),
	.col_reg_0(row3[111]),
	.col_reg_1(row3[112]),
	.col_reg_2(row3[113]),
	.col_reg_3(row3[114]),
	.col_reg_4(row3[115]),
	.col_reg_5(row3[116]),
	.col_reg_6(row3[117]),
	.col_reg_7(row3[118]),
	.col_reg_8(row3[119]),
	.col_reg_9(row3[120]),
	.col_reg_10(row3[121]),
	.col_reg_11(row3[122]),
	.col_reg_12(row3[123]),
	.col_reg_13(row3[124]),
	.col_reg_14(row3[125]),
	.col_reg_15(row3[126]),
	.col_reg_16(row3[127]),
	.col_reg_17(row3[128]),
	.col_reg_18(row3[129]),
	.col_reg_19(row3[130]),
	.col_reg_20(row3[131]),
	.col_reg_21(row3[132]),
	.col_reg_22(row3[133]),
	.col_reg_23(row3[134]),
	.col_reg_24(row3[135]),
	.col_reg_25(row3[136]),
	.col_reg_26(row3[137]),
	.col_reg_27(row3[138]),
	.col_reg_28(row3[139]),
	.col_reg_29(row3[140]),
	.col_reg_30(row3[141]),
	.col_reg_31(row3[142]),
	.col_reg_32(row3[143]),
	.col_reg_33(row3[144]),
	.col_reg_34(row3[145]),
	.col_reg_35(row3[146]),
	.col_reg_36(row3[147]),
	.col_reg_37(row3[148]),
	.col_reg_38(row3[149]),
	.col_reg_39(row3[150]),
	.col_reg_40(row3[151]),
	.col_reg_41(row3[152]),
	.col_reg_42(row3[153]),
	.col_reg_43(row3[154]),
	.col_reg_44(row3[155]),
	.col_reg_45(row3[156]),
	.col_reg_46(row3[157]),
	.col_reg_47(row3[158]),
	.col_reg_48(row3[159]),
	.col_reg_49(row3[160])
);


vga_gen_col col_row3_char4(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_28),
	.col_reg_0(row3[164]),
	.col_reg_1(row3[165]),
	.col_reg_2(row3[166]),
	.col_reg_3(row3[167]),
	.col_reg_4(row3[168]),
	.col_reg_5(row3[169]),
	.col_reg_6(row3[170]),
	.col_reg_7(row3[171]),
	.col_reg_8(row3[172]),
	.col_reg_9(row3[173]),
	.col_reg_10(row3[174]),
	.col_reg_11(row3[175]),
	.col_reg_12(row3[176]),
	.col_reg_13(row3[177]),
	.col_reg_14(row3[178]),
	.col_reg_15(row3[179]),
	.col_reg_16(row3[180]),
	.col_reg_17(row3[181]),
	.col_reg_18(row3[182]),
	.col_reg_19(row3[183]),
	.col_reg_20(row3[184]),
	.col_reg_21(row3[185]),
	.col_reg_22(row3[186]),
	.col_reg_23(row3[187]),
	.col_reg_24(row3[188]),
	.col_reg_25(row3[189]),
	.col_reg_26(row3[190]),
	.col_reg_27(row3[191]),
	.col_reg_28(row3[192]),
	.col_reg_29(row3[193]),
	.col_reg_30(row3[194]),
	.col_reg_31(row3[195]),
	.col_reg_32(row3[196]),
	.col_reg_33(row3[197]),
	.col_reg_34(row3[198]),
	.col_reg_35(row3[199]),
	.col_reg_36(row3[200]),
	.col_reg_37(row3[201]),
	.col_reg_38(row3[202]),
	.col_reg_39(row3[203]),
	.col_reg_40(row3[204]),
	.col_reg_41(row3[205]),
	.col_reg_42(row3[206]),
	.col_reg_43(row3[207]),
	.col_reg_44(row3[208]),
	.col_reg_45(row3[209]),
	.col_reg_46(row3[210]),
	.col_reg_47(row3[211]),
	.col_reg_48(row3[212]),
	.col_reg_49(row3[213])
);


vga_gen_col col_row3_char5(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_29),
	.col_reg_0(row3[217]),
	.col_reg_1(row3[218]),
	.col_reg_2(row3[219]),
	.col_reg_3(row3[220]),
	.col_reg_4(row3[221]),
	.col_reg_5(row3[222]),
	.col_reg_6(row3[223]),
	.col_reg_7(row3[224]),
	.col_reg_8(row3[225]),
	.col_reg_9(row3[226]),
	.col_reg_10(row3[227]),
	.col_reg_11(row3[228]),
	.col_reg_12(row3[229]),
	.col_reg_13(row3[230]),
	.col_reg_14(row3[231]),
	.col_reg_15(row3[232]),
	.col_reg_16(row3[233]),
	.col_reg_17(row3[234]),
	.col_reg_18(row3[235]),
	.col_reg_19(row3[236]),
	.col_reg_20(row3[237]),
	.col_reg_21(row3[238]),
	.col_reg_22(row3[239]),
	.col_reg_23(row3[240]),
	.col_reg_24(row3[241]),
	.col_reg_25(row3[242]),
	.col_reg_26(row3[243]),
	.col_reg_27(row3[244]),
	.col_reg_28(row3[245]),
	.col_reg_29(row3[246]),
	.col_reg_30(row3[247]),
	.col_reg_31(row3[248]),
	.col_reg_32(row3[249]),
	.col_reg_33(row3[250]),
	.col_reg_34(row3[251]),
	.col_reg_35(row3[252]),
	.col_reg_36(row3[253]),
	.col_reg_37(row3[254]),
	.col_reg_38(row3[255]),
	.col_reg_39(row3[256]),
	.col_reg_40(row3[257]),
	.col_reg_41(row3[258]),
	.col_reg_42(row3[259]),
	.col_reg_43(row3[260]),
	.col_reg_44(row3[261]),
	.col_reg_45(row3[262]),
	.col_reg_46(row3[263]),
	.col_reg_47(row3[264]),
	.col_reg_48(row3[265]),
	.col_reg_49(row3[266])
);


vga_gen_col col_row3_char6(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_30),
	.col_reg_0(row3[270]),
	.col_reg_1(row3[271]),
	.col_reg_2(row3[272]),
	.col_reg_3(row3[273]),
	.col_reg_4(row3[274]),
	.col_reg_5(row3[275]),
	.col_reg_6(row3[276]),
	.col_reg_7(row3[277]),
	.col_reg_8(row3[278]),
	.col_reg_9(row3[279]),
	.col_reg_10(row3[280]),
	.col_reg_11(row3[281]),
	.col_reg_12(row3[282]),
	.col_reg_13(row3[283]),
	.col_reg_14(row3[284]),
	.col_reg_15(row3[285]),
	.col_reg_16(row3[286]),
	.col_reg_17(row3[287]),
	.col_reg_18(row3[288]),
	.col_reg_19(row3[289]),
	.col_reg_20(row3[290]),
	.col_reg_21(row3[291]),
	.col_reg_22(row3[292]),
	.col_reg_23(row3[293]),
	.col_reg_24(row3[294]),
	.col_reg_25(row3[295]),
	.col_reg_26(row3[296]),
	.col_reg_27(row3[297]),
	.col_reg_28(row3[298]),
	.col_reg_29(row3[299]),
	.col_reg_30(row3[300]),
	.col_reg_31(row3[301]),
	.col_reg_32(row3[302]),
	.col_reg_33(row3[303]),
	.col_reg_34(row3[304]),
	.col_reg_35(row3[305]),
	.col_reg_36(row3[306]),
	.col_reg_37(row3[307]),
	.col_reg_38(row3[308]),
	.col_reg_39(row3[309]),
	.col_reg_40(row3[310]),
	.col_reg_41(row3[311]),
	.col_reg_42(row3[312]),
	.col_reg_43(row3[313]),
	.col_reg_44(row3[314]),
	.col_reg_45(row3[315]),
	.col_reg_46(row3[316]),
	.col_reg_47(row3[317]),
	.col_reg_48(row3[318]),
	.col_reg_49(row3[319])
);


vga_gen_col col_row3_char7(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_31),
	.col_reg_0(row3[323]),
	.col_reg_1(row3[324]),
	.col_reg_2(row3[325]),
	.col_reg_3(row3[326]),
	.col_reg_4(row3[327]),
	.col_reg_5(row3[328]),
	.col_reg_6(row3[329]),
	.col_reg_7(row3[330]),
	.col_reg_8(row3[331]),
	.col_reg_9(row3[332]),
	.col_reg_10(row3[333]),
	.col_reg_11(row3[334]),
	.col_reg_12(row3[335]),
	.col_reg_13(row3[336]),
	.col_reg_14(row3[337]),
	.col_reg_15(row3[338]),
	.col_reg_16(row3[339]),
	.col_reg_17(row3[340]),
	.col_reg_18(row3[341]),
	.col_reg_19(row3[342]),
	.col_reg_20(row3[343]),
	.col_reg_21(row3[344]),
	.col_reg_22(row3[345]),
	.col_reg_23(row3[346]),
	.col_reg_24(row3[347]),
	.col_reg_25(row3[348]),
	.col_reg_26(row3[349]),
	.col_reg_27(row3[350]),
	.col_reg_28(row3[351]),
	.col_reg_29(row3[352]),
	.col_reg_30(row3[353]),
	.col_reg_31(row3[354]),
	.col_reg_32(row3[355]),
	.col_reg_33(row3[356]),
	.col_reg_34(row3[357]),
	.col_reg_35(row3[358]),
	.col_reg_36(row3[359]),
	.col_reg_37(row3[360]),
	.col_reg_38(row3[361]),
	.col_reg_39(row3[362]),
	.col_reg_40(row3[363]),
	.col_reg_41(row3[364]),
	.col_reg_42(row3[365]),
	.col_reg_43(row3[366]),
	.col_reg_44(row3[367]),
	.col_reg_45(row3[368]),
	.col_reg_46(row3[369]),
	.col_reg_47(row3[370]),
	.col_reg_48(row3[371]),
	.col_reg_49(row3[372])
);


vga_gen_col col_row3_char8(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_32),
	.col_reg_0(row3[376]),
	.col_reg_1(row3[377]),
	.col_reg_2(row3[378]),
	.col_reg_3(row3[379]),
	.col_reg_4(row3[380]),
	.col_reg_5(row3[381]),
	.col_reg_6(row3[382]),
	.col_reg_7(row3[383]),
	.col_reg_8(row3[384]),
	.col_reg_9(row3[385]),
	.col_reg_10(row3[386]),
	.col_reg_11(row3[387]),
	.col_reg_12(row3[388]),
	.col_reg_13(row3[389]),
	.col_reg_14(row3[390]),
	.col_reg_15(row3[391]),
	.col_reg_16(row3[392]),
	.col_reg_17(row3[393]),
	.col_reg_18(row3[394]),
	.col_reg_19(row3[395]),
	.col_reg_20(row3[396]),
	.col_reg_21(row3[397]),
	.col_reg_22(row3[398]),
	.col_reg_23(row3[399]),
	.col_reg_24(row3[400]),
	.col_reg_25(row3[401]),
	.col_reg_26(row3[402]),
	.col_reg_27(row3[403]),
	.col_reg_28(row3[404]),
	.col_reg_29(row3[405]),
	.col_reg_30(row3[406]),
	.col_reg_31(row3[407]),
	.col_reg_32(row3[408]),
	.col_reg_33(row3[409]),
	.col_reg_34(row3[410]),
	.col_reg_35(row3[411]),
	.col_reg_36(row3[412]),
	.col_reg_37(row3[413]),
	.col_reg_38(row3[414]),
	.col_reg_39(row3[415]),
	.col_reg_40(row3[416]),
	.col_reg_41(row3[417]),
	.col_reg_42(row3[418]),
	.col_reg_43(row3[419]),
	.col_reg_44(row3[420]),
	.col_reg_45(row3[421]),
	.col_reg_46(row3[422]),
	.col_reg_47(row3[423]),
	.col_reg_48(row3[424]),
	.col_reg_49(row3[425])
);


vga_gen_col col_row3_char9(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_33),
	.col_reg_0(row3[429]),
	.col_reg_1(row3[430]),
	.col_reg_2(row3[431]),
	.col_reg_3(row3[432]),
	.col_reg_4(row3[433]),
	.col_reg_5(row3[434]),
	.col_reg_6(row3[435]),
	.col_reg_7(row3[436]),
	.col_reg_8(row3[437]),
	.col_reg_9(row3[438]),
	.col_reg_10(row3[439]),
	.col_reg_11(row3[440]),
	.col_reg_12(row3[441]),
	.col_reg_13(row3[442]),
	.col_reg_14(row3[443]),
	.col_reg_15(row3[444]),
	.col_reg_16(row3[445]),
	.col_reg_17(row3[446]),
	.col_reg_18(row3[447]),
	.col_reg_19(row3[448]),
	.col_reg_20(row3[449]),
	.col_reg_21(row3[450]),
	.col_reg_22(row3[451]),
	.col_reg_23(row3[452]),
	.col_reg_24(row3[453]),
	.col_reg_25(row3[454]),
	.col_reg_26(row3[455]),
	.col_reg_27(row3[456]),
	.col_reg_28(row3[457]),
	.col_reg_29(row3[458]),
	.col_reg_30(row3[459]),
	.col_reg_31(row3[460]),
	.col_reg_32(row3[461]),
	.col_reg_33(row3[462]),
	.col_reg_34(row3[463]),
	.col_reg_35(row3[464]),
	.col_reg_36(row3[465]),
	.col_reg_37(row3[466]),
	.col_reg_38(row3[467]),
	.col_reg_39(row3[468]),
	.col_reg_40(row3[469]),
	.col_reg_41(row3[470]),
	.col_reg_42(row3[471]),
	.col_reg_43(row3[472]),
	.col_reg_44(row3[473]),
	.col_reg_45(row3[474]),
	.col_reg_46(row3[475]),
	.col_reg_47(row3[476]),
	.col_reg_48(row3[477]),
	.col_reg_49(row3[478])
);


vga_gen_col col_row3_char10(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_34),
	.col_reg_0(row3[482]),
	.col_reg_1(row3[483]),
	.col_reg_2(row3[484]),
	.col_reg_3(row3[485]),
	.col_reg_4(row3[486]),
	.col_reg_5(row3[487]),
	.col_reg_6(row3[488]),
	.col_reg_7(row3[489]),
	.col_reg_8(row3[490]),
	.col_reg_9(row3[491]),
	.col_reg_10(row3[492]),
	.col_reg_11(row3[493]),
	.col_reg_12(row3[494]),
	.col_reg_13(row3[495]),
	.col_reg_14(row3[496]),
	.col_reg_15(row3[497]),
	.col_reg_16(row3[498]),
	.col_reg_17(row3[499]),
	.col_reg_18(row3[500]),
	.col_reg_19(row3[501]),
	.col_reg_20(row3[502]),
	.col_reg_21(row3[503]),
	.col_reg_22(row3[504]),
	.col_reg_23(row3[505]),
	.col_reg_24(row3[506]),
	.col_reg_25(row3[507]),
	.col_reg_26(row3[508]),
	.col_reg_27(row3[509]),
	.col_reg_28(row3[510]),
	.col_reg_29(row3[511]),
	.col_reg_30(row3[512]),
	.col_reg_31(row3[513]),
	.col_reg_32(row3[514]),
	.col_reg_33(row3[515]),
	.col_reg_34(row3[516]),
	.col_reg_35(row3[517]),
	.col_reg_36(row3[518]),
	.col_reg_37(row3[519]),
	.col_reg_38(row3[520]),
	.col_reg_39(row3[521]),
	.col_reg_40(row3[522]),
	.col_reg_41(row3[523]),
	.col_reg_42(row3[524]),
	.col_reg_43(row3[525]),
	.col_reg_44(row3[526]),
	.col_reg_45(row3[527]),
	.col_reg_46(row3[528]),
	.col_reg_47(row3[529]),
	.col_reg_48(row3[530]),
	.col_reg_49(row3[531])
);


vga_gen_col col_row3_char11(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_35),
	.col_reg_0(row3[535]),
	.col_reg_1(row3[536]),
	.col_reg_2(row3[537]),
	.col_reg_3(row3[538]),
	.col_reg_4(row3[539]),
	.col_reg_5(row3[540]),
	.col_reg_6(row3[541]),
	.col_reg_7(row3[542]),
	.col_reg_8(row3[543]),
	.col_reg_9(row3[544]),
	.col_reg_10(row3[545]),
	.col_reg_11(row3[546]),
	.col_reg_12(row3[547]),
	.col_reg_13(row3[548]),
	.col_reg_14(row3[549]),
	.col_reg_15(row3[550]),
	.col_reg_16(row3[551]),
	.col_reg_17(row3[552]),
	.col_reg_18(row3[553]),
	.col_reg_19(row3[554]),
	.col_reg_20(row3[555]),
	.col_reg_21(row3[556]),
	.col_reg_22(row3[557]),
	.col_reg_23(row3[558]),
	.col_reg_24(row3[559]),
	.col_reg_25(row3[560]),
	.col_reg_26(row3[561]),
	.col_reg_27(row3[562]),
	.col_reg_28(row3[563]),
	.col_reg_29(row3[564]),
	.col_reg_30(row3[565]),
	.col_reg_31(row3[566]),
	.col_reg_32(row3[567]),
	.col_reg_33(row3[568]),
	.col_reg_34(row3[569]),
	.col_reg_35(row3[570]),
	.col_reg_36(row3[571]),
	.col_reg_37(row3[572]),
	.col_reg_38(row3[573]),
	.col_reg_39(row3[574]),
	.col_reg_40(row3[575]),
	.col_reg_41(row3[576]),
	.col_reg_42(row3[577]),
	.col_reg_43(row3[578]),
	.col_reg_44(row3[579]),
	.col_reg_45(row3[580]),
	.col_reg_46(row3[581]),
	.col_reg_47(row3[582]),
	.col_reg_48(row3[583]),
	.col_reg_49(row3[584])
);


vga_gen_col col_row3_char12(
	.clk(clk),
	.rst_n(rst_n),
	.input_ascii(char_36),
	.col_reg_0(row3[588]),
	.col_reg_1(row3[589]),
	.col_reg_2(row3[590]),
	.col_reg_3(row3[591]),
	.col_reg_4(row3[592]),
	.col_reg_5(row3[593]),
	.col_reg_6(row3[594]),
	.col_reg_7(row3[595]),
	.col_reg_8(row3[596]),
	.col_reg_9(row3[597]),
	.col_reg_10(row3[598]),
	.col_reg_11(row3[599]),
	.col_reg_12(row3[600]),
	.col_reg_13(row3[601]),
	.col_reg_14(row3[602]),
	.col_reg_15(row3[603]),
	.col_reg_16(row3[604]),
	.col_reg_17(row3[605]),
	.col_reg_18(row3[606]),
	.col_reg_19(row3[607]),
	.col_reg_20(row3[608]),
	.col_reg_21(row3[609]),
	.col_reg_22(row3[610]),
	.col_reg_23(row3[611]),
	.col_reg_24(row3[612]),
	.col_reg_25(row3[613]),
	.col_reg_26(row3[614]),
	.col_reg_27(row3[615]),
	.col_reg_28(row3[616]),
	.col_reg_29(row3[617]),
	.col_reg_30(row3[618]),
	.col_reg_31(row3[619]),
	.col_reg_32(row3[620]),
	.col_reg_33(row3[621]),
	.col_reg_34(row3[622]),
	.col_reg_35(row3[623]),
	.col_reg_36(row3[624]),
	.col_reg_37(row3[625]),
	.col_reg_38(row3[626]),
	.col_reg_39(row3[627]),
	.col_reg_40(row3[628]),
	.col_reg_41(row3[629]),
	.col_reg_42(row3[630]),
	.col_reg_43(row3[631]),
	.col_reg_44(row3[632]),
	.col_reg_45(row3[633]),
	.col_reg_46(row3[634]),
	.col_reg_47(row3[635]),
	.col_reg_48(row3[636]),
	.col_reg_49(row3[637])
);

	always @ (posedge vga_clk or negedge rst_n)
	begin
		if (!rst_n) begin
			vga_r <= 0;
			vga_g <= 0;
			vga_b <= 0;
		end
		else 
            if (pixel_x>=LEFT_BOUND) begin // && pixel_x<=RIGHT_BOUND && pixel_y>=UP_BOUND && pixel_y<=DOWN_BOUND) begin // 如果是在显示区域
                if (pixel_y>=up_pos_row1 && pixel_y<=down_pos_row1) begin
                    if (row1[pixel_x][69-(pixel_y-up_pos_row1)]) begin
                        vga_r <= 3'b111;
                        vga_g <= 3'b111;
                        vga_b <= 3'b111;
                    end
                    else begin
                        vga_r <= 3'b000;
                        vga_g <= 3'b000;
                        vga_b <= 3'b000;
                    end
                end

                else if (pixel_y>=up_pos_row2 && pixel_y<=down_pos_row2) begin
                    if (row2[pixel_x][69-(pixel_y-up_pos_row2)]) begin
                        vga_r <= 3'b111;
                        vga_g <= 3'b111;
                        vga_b <= 3'b111;
                    end
                    else begin
                        vga_r <= 3'b000;
                        vga_g <= 3'b000;
                        vga_b <= 3'b000;
                    end
                end

                else if (pixel_y>=up_pos_row3 && pixel_y<=down_pos_row3) begin
                    if (row3[pixel_x][69-(pixel_y-up_pos_row3)]) begin
                        vga_r <= 3'b111;
                        vga_g <= 3'b111;
                        vga_b <= 3'b111;
                    end
                    else begin
                        vga_r <= 3'b000;
                        vga_g <= 3'b000;
                        vga_b <= 3'b000;
                    end
                end


                else begin
                    vga_r <= 3'b000;
                    vga_g <= 3'b000;
                    vga_b <= 3'b000;
                end
            end
            else begin
                vga_r <= 3'b000;
                vga_g <= 3'b000;
                vga_b <= 3'b000;
            end
	end

endmodule
